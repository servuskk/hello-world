library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity LAB8_voltage is

port
	(
		clk_v: in std_logic;
		rst_v: in std_logic;	
		flag: in std_logic;								--������ʾģʽ
		vin: in std_logic_vector(7 downto 0);			--ADC�õ��ģ�ͬled��ʾ�����֣��õ�ʱ����Ҫȡ��
		bcdin: in std_logic_vector(11 downto 0);
		lcdbcd: buffer std_logic_vector(19 downto 0);
-----------�����74hc595���źţ�������ʾģʽ��3.3 256��-------------------------------------
		out0: out std_logic_vector(7 downto 0);
		out1: out std_logic_vector(7 downto 0);
		out2: out std_logic_vector(7 downto 0);
		out3: out std_logic_vector(7 downto 0);
		out4: out std_logic_vector(7 downto 0);
		out5: out std_logic_vector(7 downto 0)
		
	);
end LAB8_voltage;

architecture behavior of LAB8_voltage is
	signal v_33_1: integer;
	signal v_33_2: integer;
	signal v_33_3: integer;
	signal v_33_4: integer;
	signal v_33_5: integer;
begin
	process(clk_v)
	begin
		case not vin is--ö�ٷ�yyds
			when "00000000"=> v_33_1<=0; v_33_2<=0; v_33_3<=0; v_33_4<=0; v_33_5<=0;
			when "00000001"=> v_33_1<=0; v_33_2<=0; v_33_3<=1; v_33_4<=2; v_33_5<=9;
			when "00000010"=> v_33_1<=0; v_33_2<=0; v_33_3<=2; v_33_4<=5; v_33_5<=8;
			when "00000011"=> v_33_1<=0; v_33_2<=0; v_33_3<=3; v_33_4<=8; v_33_5<=8;
			when "00000100"=> v_33_1<=0; v_33_2<=0; v_33_3<=5; v_33_4<=1; v_33_5<=7;
			when "00000101"=> v_33_1<=0; v_33_2<=0; v_33_3<=6; v_33_4<=4; v_33_5<=7;
			when "00000110"=> v_33_1<=0; v_33_2<=0; v_33_3<=7; v_33_4<=7; v_33_5<=6;
			when "00000111"=> v_33_1<=0; v_33_2<=0; v_33_3<=9; v_33_4<=0; v_33_5<=5;
			when "00001000"=> v_33_1<=0; v_33_2<=1; v_33_3<=0; v_33_4<=3; v_33_5<=5;
			when "00001001"=> v_33_1<=0; v_33_2<=1; v_33_3<=1; v_33_4<=6; v_33_5<=4;
			when "00001010"=> v_33_1<=0; v_33_2<=1; v_33_3<=2; v_33_4<=9; v_33_5<=4;
			when "00001011"=> v_33_1<=0; v_33_2<=1; v_33_3<=4; v_33_4<=2; v_33_5<=3;
			when "00001100"=> v_33_1<=0; v_33_2<=1; v_33_3<=5; v_33_4<=5; v_33_5<=2;
			when "00001101"=> v_33_1<=0; v_33_2<=1; v_33_3<=6; v_33_4<=8; v_33_5<=2;
			when "00001110"=> v_33_1<=0; v_33_2<=1; v_33_3<=8; v_33_4<=1; v_33_5<=1;
			when "00001111"=> v_33_1<=0; v_33_2<=1; v_33_3<=9; v_33_4<=4; v_33_5<=1;
			when "00010000"=> v_33_1<=0; v_33_2<=2; v_33_3<=0; v_33_4<=7; v_33_5<=0;
			when "00010001"=> v_33_1<=0; v_33_2<=2; v_33_3<=2; v_33_4<=0; v_33_5<=0;
			when "00010010"=> v_33_1<=0; v_33_2<=2; v_33_3<=3; v_33_4<=2; v_33_5<=9;
			when "00010011"=> v_33_1<=0; v_33_2<=2; v_33_3<=4; v_33_4<=5; v_33_5<=8;
			when "00010100"=> v_33_1<=0; v_33_2<=2; v_33_3<=5; v_33_4<=8; v_33_5<=8;
			when "00010101"=> v_33_1<=0; v_33_2<=2; v_33_3<=7; v_33_4<=1; v_33_5<=7;
			when "00010110"=> v_33_1<=0; v_33_2<=2; v_33_3<=8; v_33_4<=4; v_33_5<=7;
			when "00010111"=> v_33_1<=0; v_33_2<=2; v_33_3<=9; v_33_4<=7; v_33_5<=6;
			when "00011000"=> v_33_1<=0; v_33_2<=3; v_33_3<=1; v_33_4<=0; v_33_5<=5;
			when "00011001"=> v_33_1<=0; v_33_2<=3; v_33_3<=2; v_33_4<=3; v_33_5<=5;
			when "00011010"=> v_33_1<=0; v_33_2<=3; v_33_3<=3; v_33_4<=6; v_33_5<=4;
			when "00011011"=> v_33_1<=0; v_33_2<=3; v_33_3<=4; v_33_4<=9; v_33_5<=4;
			when "00011100"=> v_33_1<=0; v_33_2<=3; v_33_3<=6; v_33_4<=2; v_33_5<=3;
			when "00011101"=> v_33_1<=0; v_33_2<=3; v_33_3<=7; v_33_4<=5; v_33_5<=2;
			when "00011110"=> v_33_1<=0; v_33_2<=3; v_33_3<=8; v_33_4<=8; v_33_5<=2;
			when "00011111"=> v_33_1<=0; v_33_2<=4; v_33_3<=0; v_33_4<=1; v_33_5<=1;
			when "00100000"=> v_33_1<=0; v_33_2<=4; v_33_3<=1; v_33_4<=4; v_33_5<=1;
			when "00100001"=> v_33_1<=0; v_33_2<=4; v_33_3<=2; v_33_4<=7; v_33_5<=0;
			when "00100010"=> v_33_1<=0; v_33_2<=4; v_33_3<=4; v_33_4<=0; v_33_5<=0;
			when "00100011"=> v_33_1<=0; v_33_2<=4; v_33_3<=5; v_33_4<=2; v_33_5<=9;
			when "00100100"=> v_33_1<=0; v_33_2<=4; v_33_3<=6; v_33_4<=5; v_33_5<=8;
			when "00100101"=> v_33_1<=0; v_33_2<=4; v_33_3<=7; v_33_4<=8; v_33_5<=8;
			when "00100110"=> v_33_1<=0; v_33_2<=4; v_33_3<=9; v_33_4<=1; v_33_5<=7;
			when "00100111"=> v_33_1<=0; v_33_2<=5; v_33_3<=0; v_33_4<=4; v_33_5<=7;
			when "00101000"=> v_33_1<=0; v_33_2<=5; v_33_3<=1; v_33_4<=7; v_33_5<=6;
			when "00101001"=> v_33_1<=0; v_33_2<=5; v_33_3<=3; v_33_4<=0; v_33_5<=5;
			when "00101010"=> v_33_1<=0; v_33_2<=5; v_33_3<=4; v_33_4<=3; v_33_5<=5;
			when "00101011"=> v_33_1<=0; v_33_2<=5; v_33_3<=5; v_33_4<=6; v_33_5<=4;
			when "00101100"=> v_33_1<=0; v_33_2<=5; v_33_3<=6; v_33_4<=9; v_33_5<=4;
			when "00101101"=> v_33_1<=0; v_33_2<=5; v_33_3<=8; v_33_4<=2; v_33_5<=3;
			when "00101110"=> v_33_1<=0; v_33_2<=5; v_33_3<=9; v_33_4<=5; v_33_5<=2;
			when "00101111"=> v_33_1<=0; v_33_2<=6; v_33_3<=0; v_33_4<=8; v_33_5<=2;
			when "00110000"=> v_33_1<=0; v_33_2<=6; v_33_3<=2; v_33_4<=1; v_33_5<=1;
			when "00110001"=> v_33_1<=0; v_33_2<=6; v_33_3<=3; v_33_4<=4; v_33_5<=1;
			when "00110010"=> v_33_1<=0; v_33_2<=6; v_33_3<=4; v_33_4<=7; v_33_5<=0;
			when "00110011"=> v_33_1<=0; v_33_2<=6; v_33_3<=6; v_33_4<=0; v_33_5<=0;
			when "00110100"=> v_33_1<=0; v_33_2<=6; v_33_3<=7; v_33_4<=2; v_33_5<=9;
			when "00110101"=> v_33_1<=0; v_33_2<=6; v_33_3<=8; v_33_4<=5; v_33_5<=8;
			when "00110110"=> v_33_1<=0; v_33_2<=6; v_33_3<=9; v_33_4<=8; v_33_5<=8;
			when "00110111"=> v_33_1<=0; v_33_2<=7; v_33_3<=1; v_33_4<=1; v_33_5<=7;
			when "00111000"=> v_33_1<=0; v_33_2<=7; v_33_3<=2; v_33_4<=4; v_33_5<=7;
			when "00111001"=> v_33_1<=0; v_33_2<=7; v_33_3<=3; v_33_4<=7; v_33_5<=6;
			when "00111010"=> v_33_1<=0; v_33_2<=7; v_33_3<=5; v_33_4<=0; v_33_5<=5;
			when "00111011"=> v_33_1<=0; v_33_2<=7; v_33_3<=6; v_33_4<=3; v_33_5<=5;
			when "00111100"=> v_33_1<=0; v_33_2<=7; v_33_3<=7; v_33_4<=6; v_33_5<=4;
			when "00111101"=> v_33_1<=0; v_33_2<=7; v_33_3<=8; v_33_4<=9; v_33_5<=4;
			when "00111110"=> v_33_1<=0; v_33_2<=8; v_33_3<=0; v_33_4<=2; v_33_5<=3;
			when "00111111"=> v_33_1<=0; v_33_2<=8; v_33_3<=1; v_33_4<=5; v_33_5<=2;
			when "01000000"=> v_33_1<=0; v_33_2<=8; v_33_3<=2; v_33_4<=8; v_33_5<=2;
			when "01000001"=> v_33_1<=0; v_33_2<=8; v_33_3<=4; v_33_4<=1; v_33_5<=1;
			when "01000010"=> v_33_1<=0; v_33_2<=8; v_33_3<=5; v_33_4<=4; v_33_5<=1;
			when "01000011"=> v_33_1<=0; v_33_2<=8; v_33_3<=6; v_33_4<=7; v_33_5<=0;
			when "01000100"=> v_33_1<=0; v_33_2<=8; v_33_3<=8; v_33_4<=0; v_33_5<=0;
			when "01000101"=> v_33_1<=0; v_33_2<=8; v_33_3<=9; v_33_4<=2; v_33_5<=9;
			when "01000110"=> v_33_1<=0; v_33_2<=9; v_33_3<=0; v_33_4<=5; v_33_5<=8;
			when "01000111"=> v_33_1<=0; v_33_2<=9; v_33_3<=1; v_33_4<=8; v_33_5<=8;
			when "01001000"=> v_33_1<=0; v_33_2<=9; v_33_3<=3; v_33_4<=1; v_33_5<=7;
			when "01001001"=> v_33_1<=0; v_33_2<=9; v_33_3<=4; v_33_4<=4; v_33_5<=7;
			when "01001010"=> v_33_1<=0; v_33_2<=9; v_33_3<=5; v_33_4<=7; v_33_5<=6;
			when "01001011"=> v_33_1<=0; v_33_2<=9; v_33_3<=7; v_33_4<=0; v_33_5<=5;
			when "01001100"=> v_33_1<=0; v_33_2<=9; v_33_3<=8; v_33_4<=3; v_33_5<=5;
			when "01001101"=> v_33_1<=0; v_33_2<=9; v_33_3<=9; v_33_4<=6; v_33_5<=4;
			when "01001110"=> v_33_1<=1; v_33_2<=0; v_33_3<=0; v_33_4<=9; v_33_5<=4;
			when "01001111"=> v_33_1<=1; v_33_2<=0; v_33_3<=2; v_33_4<=2; v_33_5<=3;
			when "01010000"=> v_33_1<=1; v_33_2<=0; v_33_3<=3; v_33_4<=5; v_33_5<=2;
			when "01010001"=> v_33_1<=1; v_33_2<=0; v_33_3<=4; v_33_4<=8; v_33_5<=2;
			when "01010010"=> v_33_1<=1; v_33_2<=0; v_33_3<=6; v_33_4<=1; v_33_5<=1;
			when "01010011"=> v_33_1<=1; v_33_2<=0; v_33_3<=7; v_33_4<=4; v_33_5<=1;
			when "01010100"=> v_33_1<=1; v_33_2<=0; v_33_3<=8; v_33_4<=7; v_33_5<=0;
			when "01010101"=> v_33_1<=1; v_33_2<=1; v_33_3<=0; v_33_4<=0; v_33_5<=0;
			when "01010110"=> v_33_1<=1; v_33_2<=1; v_33_3<=1; v_33_4<=2; v_33_5<=9;
			when "01010111"=> v_33_1<=1; v_33_2<=1; v_33_3<=2; v_33_4<=5; v_33_5<=8;
			when "01011000"=> v_33_1<=1; v_33_2<=1; v_33_3<=3; v_33_4<=8; v_33_5<=8;
			when "01011001"=> v_33_1<=1; v_33_2<=1; v_33_3<=5; v_33_4<=1; v_33_5<=7;
			when "01011010"=> v_33_1<=1; v_33_2<=1; v_33_3<=6; v_33_4<=4; v_33_5<=7;
			when "01011011"=> v_33_1<=1; v_33_2<=1; v_33_3<=7; v_33_4<=7; v_33_5<=6;
			when "01011100"=> v_33_1<=1; v_33_2<=1; v_33_3<=9; v_33_4<=0; v_33_5<=5;
			when "01011101"=> v_33_1<=1; v_33_2<=2; v_33_3<=0; v_33_4<=3; v_33_5<=5;
			when "01011110"=> v_33_1<=1; v_33_2<=2; v_33_3<=1; v_33_4<=6; v_33_5<=4;
			when "01011111"=> v_33_1<=1; v_33_2<=2; v_33_3<=2; v_33_4<=9; v_33_5<=4;
			when "01100000"=> v_33_1<=1; v_33_2<=2; v_33_3<=4; v_33_4<=2; v_33_5<=3;
			when "01100001"=> v_33_1<=1; v_33_2<=2; v_33_3<=5; v_33_4<=5; v_33_5<=2;
			when "01100010"=> v_33_1<=1; v_33_2<=2; v_33_3<=6; v_33_4<=8; v_33_5<=2;
			when "01100011"=> v_33_1<=1; v_33_2<=2; v_33_3<=8; v_33_4<=1; v_33_5<=1;
			when "01100100"=> v_33_1<=1; v_33_2<=2; v_33_3<=9; v_33_4<=4; v_33_5<=1;
			when "01100101"=> v_33_1<=1; v_33_2<=3; v_33_3<=0; v_33_4<=7; v_33_5<=0;
			when "01100110"=> v_33_1<=1; v_33_2<=3; v_33_3<=2; v_33_4<=0; v_33_5<=0;
			when "01100111"=> v_33_1<=1; v_33_2<=3; v_33_3<=3; v_33_4<=2; v_33_5<=9;
			when "01101000"=> v_33_1<=1; v_33_2<=3; v_33_3<=4; v_33_4<=5; v_33_5<=8;
			when "01101001"=> v_33_1<=1; v_33_2<=3; v_33_3<=5; v_33_4<=8; v_33_5<=8;
			when "01101010"=> v_33_1<=1; v_33_2<=3; v_33_3<=7; v_33_4<=1; v_33_5<=7;
			when "01101011"=> v_33_1<=1; v_33_2<=3; v_33_3<=8; v_33_4<=4; v_33_5<=7;
			when "01101100"=> v_33_1<=1; v_33_2<=3; v_33_3<=9; v_33_4<=7; v_33_5<=6;
			when "01101101"=> v_33_1<=1; v_33_2<=4; v_33_3<=1; v_33_4<=0; v_33_5<=5;
			when "01101110"=> v_33_1<=1; v_33_2<=4; v_33_3<=2; v_33_4<=3; v_33_5<=5;
			when "01101111"=> v_33_1<=1; v_33_2<=4; v_33_3<=3; v_33_4<=6; v_33_5<=4;
			when "01110000"=> v_33_1<=1; v_33_2<=4; v_33_3<=4; v_33_4<=9; v_33_5<=4;
			when "01110001"=> v_33_1<=1; v_33_2<=4; v_33_3<=6; v_33_4<=2; v_33_5<=3;
			when "01110010"=> v_33_1<=1; v_33_2<=4; v_33_3<=7; v_33_4<=5; v_33_5<=2;
			when "01110011"=> v_33_1<=1; v_33_2<=4; v_33_3<=8; v_33_4<=8; v_33_5<=2;
			when "01110100"=> v_33_1<=1; v_33_2<=5; v_33_3<=0; v_33_4<=1; v_33_5<=1;
			when "01110101"=> v_33_1<=1; v_33_2<=5; v_33_3<=1; v_33_4<=4; v_33_5<=1;
			when "01110110"=> v_33_1<=1; v_33_2<=5; v_33_3<=2; v_33_4<=7; v_33_5<=0;
			when "01110111"=> v_33_1<=1; v_33_2<=5; v_33_3<=4; v_33_4<=0; v_33_5<=0;
			when "01111000"=> v_33_1<=1; v_33_2<=5; v_33_3<=5; v_33_4<=2; v_33_5<=9;
			when "01111001"=> v_33_1<=1; v_33_2<=5; v_33_3<=6; v_33_4<=5; v_33_5<=8;
			when "01111010"=> v_33_1<=1; v_33_2<=5; v_33_3<=7; v_33_4<=8; v_33_5<=8;
			when "01111011"=> v_33_1<=1; v_33_2<=5; v_33_3<=9; v_33_4<=1; v_33_5<=7;
			when "01111100"=> v_33_1<=1; v_33_2<=6; v_33_3<=0; v_33_4<=4; v_33_5<=7;
			when "01111101"=> v_33_1<=1; v_33_2<=6; v_33_3<=1; v_33_4<=7; v_33_5<=6;
			when "01111110"=> v_33_1<=1; v_33_2<=6; v_33_3<=3; v_33_4<=0; v_33_5<=5;
			when "01111111"=> v_33_1<=1; v_33_2<=6; v_33_3<=4; v_33_4<=3; v_33_5<=5;
			when "10000000"=> v_33_1<=1; v_33_2<=6; v_33_3<=5; v_33_4<=6; v_33_5<=4;
			when "10000001"=> v_33_1<=1; v_33_2<=6; v_33_3<=6; v_33_4<=9; v_33_5<=4;
			when "10000010"=> v_33_1<=1; v_33_2<=6; v_33_3<=8; v_33_4<=2; v_33_5<=3;
			when "10000011"=> v_33_1<=1; v_33_2<=6; v_33_3<=9; v_33_4<=5; v_33_5<=2;
			when "10000100"=> v_33_1<=1; v_33_2<=7; v_33_3<=0; v_33_4<=8; v_33_5<=2;
			when "10000101"=> v_33_1<=1; v_33_2<=7; v_33_3<=2; v_33_4<=1; v_33_5<=1;
			when "10000110"=> v_33_1<=1; v_33_2<=7; v_33_3<=3; v_33_4<=4; v_33_5<=1;
			when "10000111"=> v_33_1<=1; v_33_2<=7; v_33_3<=4; v_33_4<=7; v_33_5<=0;
			when "10001000"=> v_33_1<=1; v_33_2<=7; v_33_3<=6; v_33_4<=0; v_33_5<=0;
			when "10001001"=> v_33_1<=1; v_33_2<=7; v_33_3<=7; v_33_4<=2; v_33_5<=9;
			when "10001010"=> v_33_1<=1; v_33_2<=7; v_33_3<=8; v_33_4<=5; v_33_5<=8;
			when "10001011"=> v_33_1<=1; v_33_2<=7; v_33_3<=9; v_33_4<=8; v_33_5<=8;
			when "10001100"=> v_33_1<=1; v_33_2<=8; v_33_3<=1; v_33_4<=1; v_33_5<=7;
			when "10001101"=> v_33_1<=1; v_33_2<=8; v_33_3<=2; v_33_4<=4; v_33_5<=7;
			when "10001110"=> v_33_1<=1; v_33_2<=8; v_33_3<=3; v_33_4<=7; v_33_5<=6;
			when "10001111"=> v_33_1<=1; v_33_2<=8; v_33_3<=5; v_33_4<=0; v_33_5<=5;
			when "10010000"=> v_33_1<=1; v_33_2<=8; v_33_3<=6; v_33_4<=3; v_33_5<=5;
			when "10010001"=> v_33_1<=1; v_33_2<=8; v_33_3<=7; v_33_4<=6; v_33_5<=4;
			when "10010010"=> v_33_1<=1; v_33_2<=8; v_33_3<=8; v_33_4<=9; v_33_5<=4;
			when "10010011"=> v_33_1<=1; v_33_2<=9; v_33_3<=0; v_33_4<=2; v_33_5<=3;
			when "10010100"=> v_33_1<=1; v_33_2<=9; v_33_3<=1; v_33_4<=5; v_33_5<=2;
			when "10010101"=> v_33_1<=1; v_33_2<=9; v_33_3<=2; v_33_4<=8; v_33_5<=2;
			when "10010110"=> v_33_1<=1; v_33_2<=9; v_33_3<=4; v_33_4<=1; v_33_5<=1;
			when "10010111"=> v_33_1<=1; v_33_2<=9; v_33_3<=5; v_33_4<=4; v_33_5<=1;
			when "10011000"=> v_33_1<=1; v_33_2<=9; v_33_3<=6; v_33_4<=7; v_33_5<=0;
			when "10011001"=> v_33_1<=1; v_33_2<=9; v_33_3<=8; v_33_4<=0; v_33_5<=0;
			when "10011010"=> v_33_1<=1; v_33_2<=9; v_33_3<=9; v_33_4<=2; v_33_5<=9;
			when "10011011"=> v_33_1<=2; v_33_2<=0; v_33_3<=0; v_33_4<=5; v_33_5<=8;
			when "10011100"=> v_33_1<=2; v_33_2<=0; v_33_3<=1; v_33_4<=8; v_33_5<=8;
			when "10011101"=> v_33_1<=2; v_33_2<=0; v_33_3<=3; v_33_4<=1; v_33_5<=7;
			when "10011110"=> v_33_1<=2; v_33_2<=0; v_33_3<=4; v_33_4<=4; v_33_5<=7;
			when "10011111"=> v_33_1<=2; v_33_2<=0; v_33_3<=5; v_33_4<=7; v_33_5<=6;
			when "10100000"=> v_33_1<=2; v_33_2<=0; v_33_3<=7; v_33_4<=0; v_33_5<=5;
			when "10100001"=> v_33_1<=2; v_33_2<=0; v_33_3<=8; v_33_4<=3; v_33_5<=5;
			when "10100010"=> v_33_1<=2; v_33_2<=0; v_33_3<=9; v_33_4<=6; v_33_5<=4;
			when "10100011"=> v_33_1<=2; v_33_2<=1; v_33_3<=0; v_33_4<=9; v_33_5<=4;
			when "10100100"=> v_33_1<=2; v_33_2<=1; v_33_3<=2; v_33_4<=2; v_33_5<=3;
			when "10100101"=> v_33_1<=2; v_33_2<=1; v_33_3<=3; v_33_4<=5; v_33_5<=2;
			when "10100110"=> v_33_1<=2; v_33_2<=1; v_33_3<=4; v_33_4<=8; v_33_5<=2;
			when "10100111"=> v_33_1<=2; v_33_2<=1; v_33_3<=6; v_33_4<=1; v_33_5<=1;
			when "10101000"=> v_33_1<=2; v_33_2<=1; v_33_3<=7; v_33_4<=4; v_33_5<=1;
			when "10101001"=> v_33_1<=2; v_33_2<=1; v_33_3<=8; v_33_4<=7; v_33_5<=0;
			when "10101010"=> v_33_1<=2; v_33_2<=2; v_33_3<=0; v_33_4<=0; v_33_5<=0;
			when "10101011"=> v_33_1<=2; v_33_2<=2; v_33_3<=1; v_33_4<=2; v_33_5<=9;
			when "10101100"=> v_33_1<=2; v_33_2<=2; v_33_3<=2; v_33_4<=5; v_33_5<=8;
			when "10101101"=> v_33_1<=2; v_33_2<=2; v_33_3<=3; v_33_4<=8; v_33_5<=8;
			when "10101110"=> v_33_1<=2; v_33_2<=2; v_33_3<=5; v_33_4<=1; v_33_5<=7;
			when "10101111"=> v_33_1<=2; v_33_2<=2; v_33_3<=6; v_33_4<=4; v_33_5<=7;
			when "10110000"=> v_33_1<=2; v_33_2<=2; v_33_3<=7; v_33_4<=7; v_33_5<=6;
			when "10110001"=> v_33_1<=2; v_33_2<=2; v_33_3<=9; v_33_4<=0; v_33_5<=5;
			when "10110010"=> v_33_1<=2; v_33_2<=3; v_33_3<=0; v_33_4<=3; v_33_5<=5;
			when "10110011"=> v_33_1<=2; v_33_2<=3; v_33_3<=1; v_33_4<=6; v_33_5<=4;
			when "10110100"=> v_33_1<=2; v_33_2<=3; v_33_3<=2; v_33_4<=9; v_33_5<=4;
			when "10110101"=> v_33_1<=2; v_33_2<=3; v_33_3<=4; v_33_4<=2; v_33_5<=3;
			when "10110110"=> v_33_1<=2; v_33_2<=3; v_33_3<=5; v_33_4<=5; v_33_5<=2;
			when "10110111"=> v_33_1<=2; v_33_2<=3; v_33_3<=6; v_33_4<=8; v_33_5<=2;
			when "10111000"=> v_33_1<=2; v_33_2<=3; v_33_3<=8; v_33_4<=1; v_33_5<=1;
			when "10111001"=> v_33_1<=2; v_33_2<=3; v_33_3<=9; v_33_4<=4; v_33_5<=1;
			when "10111010"=> v_33_1<=2; v_33_2<=4; v_33_3<=0; v_33_4<=7; v_33_5<=0;
			when "10111011"=> v_33_1<=2; v_33_2<=4; v_33_3<=2; v_33_4<=0; v_33_5<=0;
			when "10111100"=> v_33_1<=2; v_33_2<=4; v_33_3<=3; v_33_4<=2; v_33_5<=9;
			when "10111101"=> v_33_1<=2; v_33_2<=4; v_33_3<=4; v_33_4<=5; v_33_5<=8;
			when "10111110"=> v_33_1<=2; v_33_2<=4; v_33_3<=5; v_33_4<=8; v_33_5<=8;
			when "10111111"=> v_33_1<=2; v_33_2<=4; v_33_3<=7; v_33_4<=1; v_33_5<=7;
			when "11000000"=> v_33_1<=2; v_33_2<=4; v_33_3<=8; v_33_4<=4; v_33_5<=7;
			when "11000001"=> v_33_1<=2; v_33_2<=4; v_33_3<=9; v_33_4<=7; v_33_5<=6;
			when "11000010"=> v_33_1<=2; v_33_2<=5; v_33_3<=1; v_33_4<=0; v_33_5<=5;
			when "11000011"=> v_33_1<=2; v_33_2<=5; v_33_3<=2; v_33_4<=3; v_33_5<=5;
			when "11000100"=> v_33_1<=2; v_33_2<=5; v_33_3<=3; v_33_4<=6; v_33_5<=4;
			when "11000101"=> v_33_1<=2; v_33_2<=5; v_33_3<=4; v_33_4<=9; v_33_5<=4;
			when "11000110"=> v_33_1<=2; v_33_2<=5; v_33_3<=6; v_33_4<=2; v_33_5<=3;
			when "11000111"=> v_33_1<=2; v_33_2<=5; v_33_3<=7; v_33_4<=5; v_33_5<=2;
			when "11001000"=> v_33_1<=2; v_33_2<=5; v_33_3<=8; v_33_4<=8; v_33_5<=2;
			when "11001001"=> v_33_1<=2; v_33_2<=6; v_33_3<=0; v_33_4<=1; v_33_5<=1;
			when "11001010"=> v_33_1<=2; v_33_2<=6; v_33_3<=1; v_33_4<=4; v_33_5<=1;
			when "11001011"=> v_33_1<=2; v_33_2<=6; v_33_3<=2; v_33_4<=7; v_33_5<=0;
			when "11001100"=> v_33_1<=2; v_33_2<=6; v_33_3<=4; v_33_4<=0; v_33_5<=0;
			when "11001101"=> v_33_1<=2; v_33_2<=6; v_33_3<=5; v_33_4<=2; v_33_5<=9;
			when "11001110"=> v_33_1<=2; v_33_2<=6; v_33_3<=6; v_33_4<=5; v_33_5<=8;
			when "11001111"=> v_33_1<=2; v_33_2<=6; v_33_3<=7; v_33_4<=8; v_33_5<=8;
			when "11010000"=> v_33_1<=2; v_33_2<=6; v_33_3<=9; v_33_4<=1; v_33_5<=7;
			when "11010001"=> v_33_1<=2; v_33_2<=7; v_33_3<=0; v_33_4<=4; v_33_5<=7;
			when "11010010"=> v_33_1<=2; v_33_2<=7; v_33_3<=1; v_33_4<=7; v_33_5<=6;
			when "11010011"=> v_33_1<=2; v_33_2<=7; v_33_3<=3; v_33_4<=0; v_33_5<=5;
			when "11010100"=> v_33_1<=2; v_33_2<=7; v_33_3<=4; v_33_4<=3; v_33_5<=5;
			when "11010101"=> v_33_1<=2; v_33_2<=7; v_33_3<=5; v_33_4<=6; v_33_5<=4;
			when "11010110"=> v_33_1<=2; v_33_2<=7; v_33_3<=6; v_33_4<=9; v_33_5<=4;
			when "11010111"=> v_33_1<=2; v_33_2<=7; v_33_3<=8; v_33_4<=2; v_33_5<=3;
			when "11011000"=> v_33_1<=2; v_33_2<=7; v_33_3<=9; v_33_4<=5; v_33_5<=2;
			when "11011001"=> v_33_1<=2; v_33_2<=8; v_33_3<=0; v_33_4<=8; v_33_5<=2;
			when "11011010"=> v_33_1<=2; v_33_2<=8; v_33_3<=2; v_33_4<=1; v_33_5<=1;
			when "11011011"=> v_33_1<=2; v_33_2<=8; v_33_3<=3; v_33_4<=4; v_33_5<=1;
			when "11011100"=> v_33_1<=2; v_33_2<=8; v_33_3<=4; v_33_4<=7; v_33_5<=0;
			when "11011101"=> v_33_1<=2; v_33_2<=8; v_33_3<=6; v_33_4<=0; v_33_5<=0;
			when "11011110"=> v_33_1<=2; v_33_2<=8; v_33_3<=7; v_33_4<=2; v_33_5<=9;
			when "11011111"=> v_33_1<=2; v_33_2<=8; v_33_3<=8; v_33_4<=5; v_33_5<=8;
			when "11100000"=> v_33_1<=2; v_33_2<=8; v_33_3<=9; v_33_4<=8; v_33_5<=8;
			when "11100001"=> v_33_1<=2; v_33_2<=9; v_33_3<=1; v_33_4<=1; v_33_5<=7;
			when "11100010"=> v_33_1<=2; v_33_2<=9; v_33_3<=2; v_33_4<=4; v_33_5<=7;
			when "11100011"=> v_33_1<=2; v_33_2<=9; v_33_3<=3; v_33_4<=7; v_33_5<=6;
			when "11100100"=> v_33_1<=2; v_33_2<=9; v_33_3<=5; v_33_4<=0; v_33_5<=5;
			when "11100101"=> v_33_1<=2; v_33_2<=9; v_33_3<=6; v_33_4<=3; v_33_5<=5;
			when "11100110"=> v_33_1<=2; v_33_2<=9; v_33_3<=7; v_33_4<=6; v_33_5<=4;
			when "11100111"=> v_33_1<=2; v_33_2<=9; v_33_3<=8; v_33_4<=9; v_33_5<=4;
			when "11101000"=> v_33_1<=3; v_33_2<=0; v_33_3<=0; v_33_4<=2; v_33_5<=3;
			when "11101001"=> v_33_1<=3; v_33_2<=0; v_33_3<=1; v_33_4<=5; v_33_5<=2;
			when "11101010"=> v_33_1<=3; v_33_2<=0; v_33_3<=2; v_33_4<=8; v_33_5<=2;
			when "11101011"=> v_33_1<=3; v_33_2<=0; v_33_3<=4; v_33_4<=1; v_33_5<=1;
			when "11101100"=> v_33_1<=3; v_33_2<=0; v_33_3<=5; v_33_4<=4; v_33_5<=1;
			when "11101101"=> v_33_1<=3; v_33_2<=0; v_33_3<=6; v_33_4<=7; v_33_5<=0;
			when "11101110"=> v_33_1<=3; v_33_2<=0; v_33_3<=8; v_33_4<=0; v_33_5<=0;
			when "11101111"=> v_33_1<=3; v_33_2<=0; v_33_3<=9; v_33_4<=2; v_33_5<=9;
			when "11110000"=> v_33_1<=3; v_33_2<=1; v_33_3<=0; v_33_4<=5; v_33_5<=8;
			when "11110001"=> v_33_1<=3; v_33_2<=1; v_33_3<=1; v_33_4<=8; v_33_5<=8;
			when "11110010"=> v_33_1<=3; v_33_2<=1; v_33_3<=3; v_33_4<=1; v_33_5<=7;
			when "11110011"=> v_33_1<=3; v_33_2<=1; v_33_3<=4; v_33_4<=4; v_33_5<=7;
			when "11110100"=> v_33_1<=3; v_33_2<=1; v_33_3<=5; v_33_4<=7; v_33_5<=6;
			when "11110101"=> v_33_1<=3; v_33_2<=1; v_33_3<=7; v_33_4<=0; v_33_5<=5;
			when "11110110"=> v_33_1<=3; v_33_2<=1; v_33_3<=8; v_33_4<=3; v_33_5<=5;
			when "11110111"=> v_33_1<=3; v_33_2<=1; v_33_3<=9; v_33_4<=6; v_33_5<=4;
			when "11111000"=> v_33_1<=3; v_33_2<=2; v_33_3<=0; v_33_4<=9; v_33_5<=4;
			when "11111001"=> v_33_1<=3; v_33_2<=2; v_33_3<=2; v_33_4<=2; v_33_5<=3;
			when "11111010"=> v_33_1<=3; v_33_2<=2; v_33_3<=3; v_33_4<=5; v_33_5<=2;
			when "11111011"=> v_33_1<=3; v_33_2<=2; v_33_3<=4; v_33_4<=8; v_33_5<=2;
			when "11111100"=> v_33_1<=3; v_33_2<=2; v_33_3<=6; v_33_4<=1; v_33_5<=1;
			when "11111101"=> v_33_1<=3; v_33_2<=2; v_33_3<=7; v_33_4<=4; v_33_5<=1;
			when "11111110"=> v_33_1<=3; v_33_2<=2; v_33_3<=8; v_33_4<=7; v_33_5<=0;
			when "11111111"=> v_33_1<=3; v_33_2<=3; v_33_3<=0; v_33_4<=0; v_33_5<=0;
			when others=> v_33_1<=0; v_33_2<=0; v_33_3<=0; v_33_4<=0; v_33_5<=0;
		end case;
	end process;
		
	process(clk_v)
		variable lcd_bcd:std_logic_vector(19 downto 0):="00000000000000000000";
	begin

			case v_33_1 is
				when 0 =>  lcd_bcd(19 downto 16):="0000";
				when 1 =>  lcd_bcd(19 downto 16):="0001";
				when 2 =>  lcd_bcd(19 downto 16):="0010";
				when 3 =>  lcd_bcd(19 downto 16):="0011";
				when 4 =>  lcd_bcd(19 downto 16):="0100";
				when 5 =>  lcd_bcd(19 downto 16):="0101";
				when 6 =>  lcd_bcd(19 downto 16):="0110";
				when 7 =>  lcd_bcd(19 downto 16):="0111";
				when 8 =>  lcd_bcd(19 downto 16):="1000";
				when 9 =>  lcd_bcd(19 downto 16):="1001";
				when others=> lcd_bcd(19 downto 16):="0000";
			end case;
			case v_33_2 is
				when 0 =>  lcd_bcd(15 downto 12):="0000";
				when 1 =>  lcd_bcd(15 downto 12):="0001";
				when 2 =>  lcd_bcd(15 downto 12):="0010";
				when 3 =>  lcd_bcd(15 downto 12):="0011";
				when 4 =>  lcd_bcd(15 downto 12):="0100";
				when 5 =>  lcd_bcd(15 downto 12):="0101";
				when 6 =>  lcd_bcd(15 downto 12):="0110";
				when 7 =>  lcd_bcd(15 downto 12):="0111";
				when 8 =>  lcd_bcd(15 downto 12):="1000";
				when 9 =>  lcd_bcd(15 downto 12):="1001";
				when others=> lcd_bcd(15 downto 12):="0000";
			end case;
			case v_33_3 is
				when 0 =>  lcd_bcd(11 downto 8):="0000";
				when 1 =>  lcd_bcd(11 downto 8):="0001";
				when 2 =>  lcd_bcd(11 downto 8):="0010";
				when 3 =>  lcd_bcd(11 downto 8):="0011";
				when 4 =>  lcd_bcd(11 downto 8):="0100";
				when 5 =>  lcd_bcd(11 downto 8):="0101";
				when 6 =>  lcd_bcd(11 downto 8):="0110";
				when 7 =>  lcd_bcd(11 downto 8):="0111";
				when 8 =>  lcd_bcd(11 downto 8):="1000";
				when 9 =>  lcd_bcd(11 downto 8):="1001";
				when others=> lcd_bcd(11 downto 8):="0000";
			end case;
			case v_33_4 is
				when 0 =>  lcd_bcd(7 downto 4):="0000";
				when 1 =>  lcd_bcd(7 downto 4):="0001";
				when 2 =>  lcd_bcd(7 downto 4):="0010";
				when 3 =>  lcd_bcd(7 downto 4):="0011";
				when 4 =>  lcd_bcd(7 downto 4):="0100";
				when 5 =>  lcd_bcd(7 downto 4):="0101";
				when 6 =>  lcd_bcd(7 downto 4):="0110";
				when 7 =>  lcd_bcd(7 downto 4):="0111";
				when 8 =>  lcd_bcd(7 downto 4):="1000";
				when 9 =>  lcd_bcd(7 downto 4):="1001";
				when others=> lcd_bcd(7 downto 4):="0000";
			end case;
			case v_33_5 is
				when 0 =>  lcd_bcd(3 downto 0):="0000";
				when 1 =>  lcd_bcd(3 downto 0):="0001";
				when 2 =>  lcd_bcd(3 downto 0):="0010";
				when 3 =>  lcd_bcd(3 downto 0):="0011";
				when 4 =>  lcd_bcd(3 downto 0):="0100";
				when 5 =>  lcd_bcd(3 downto 0):="0101";
				when 6 =>  lcd_bcd(3 downto 0):="0110";
				when 7 =>  lcd_bcd(3 downto 0):="0111";
				when 8 =>  lcd_bcd(3 downto 0):="1000";
				when 9 =>  lcd_bcd(3 downto 0):="1001";
				when others=> lcd_bcd(3 downto 0):="0000";
			end case;

		lcdbcd<=lcd_bcd;

		out0<="00000000";
------------------------------����ģʽ��ʾ----------------------------------------
		if  flag='1' then
			case v_33_1 is
				when 0 => out1<="11111101";
				when 1 => out1<="01100001";
				when 2 => out1<="11011011"; 
				when 3 => out1<="11110011";
				when 4 => out1<="01100111"; 
				when 5 => out1<="10110111";
				when 6 => out1<="10111111";
				when 7 => out1<="11100001"; 
				when 8 => out1<="11111111";
				when 9 => out1<="11110111";
				when others=>out1<="11111100";
			end case;
			case v_33_2 is
				when 0 => out2<="11111100";
				when 1 => out2<="01100000";
				when 2 => out2<="11011010"; 
				when 3 => out2<="11110010";
				when 4 => out2<="01100110"; 
				when 5 => out2<="10110110";
				when 6 => out2<="10111110";
				when 7 => out2<="11100000"; 
				when 8 => out2<="11111110";
				when 9 => out2<="11110110";
				when others=>out2<="11111100";
			end case;	
			case v_33_3 is
				when 0 => out3<="11111100";
				when 1 => out3<="01100000";
				when 2 => out3<="11011010"; 
				when 3 => out3<="11110010";
				when 4 => out3<="01100110"; 
				when 5 => out3<="10110110";
				when 6 => out3<="10111110";
				when 7 => out3<="11100000"; 
				when 8 => out3<="11111110";
				when 9 => out3<="11110110";
				when others=>out3<="11111100";
			end case;
			case v_33_4 is
				when 0 => out4<="11111100";
				when 1 => out4<="01100000";
				when 2 => out4<="11011010"; 
				when 3 => out4<="11110010";
				when 4 => out4<="01100110"; 
				when 5 => out4<="10110110";
				when 6 => out4<="10111110";
				when 7 => out4<="11100000"; 
				when 8 => out4<="11111110";
				when 9 => out4<="11110110";
				when others=>out4<="11111100";
			end case;
			case v_33_5 is
				when 0 => out5<="11111100";
				when 1 => out5<="01100000";
				when 2 => out5<="11011010"; 
				when 3 => out5<="11110010";
				when 4 => out5<="01100110"; 
				when 5 => out5<="10110110";
				when 6 => out5<="10111110";
				when 7 => out5<="11100000"; 
				when 8 => out5<="11111110";
				when 9 => out5<="11110110";
				when others=>out5<="11111100";
			end case;
		else 
			if flag='0' then----һ��Ҫ�ټ�һ��if����֪��Ϊʲô
				out1<="00000000";
				out2<="00000000";
				case bcdin(3 downto 0) is
					when "0000" => out5<= "11111100";
					when "0001" => out5<= "01100000";
					when "0010" => out5<= "11011010"; 
					when "0011" => out5<= "11110010"; 
					when "0100" => out5<= "01100110"; 
					when "0101" => out5<= "10110110";
					when "0110" => out5<= "10111110";
					when "0111" => out5<= "11100000"; 
					when "1000" => out5<= "11111110";
					when "1001" => out5<= "11110110";
					when others =>out5<= "01100000";
				end case;
				case bcdin(7 downto 4) is
					when "0000" => out4<= "11111100";
					when "0001" => out4<= "01100000";
					when "0010" => out4<= "11011010"; 
					when "0011" => out4<= "11110010"; 
					when "0100" => out4<= "01100110"; 
					when "0101" => out4<= "10110110";
					when "0110" => out4<= "10111110";
					when "0111" => out4<= "11100000"; 
					when "1000" => out4<= "11111110";
					when "1001" => out4<= "11110110";
					when others =>out4<= "01100000";
				end case;
				case bcdin(11 downto 8) is
					when "0000" => out3<= "11111100";
					when "0001" => out3<= "01100000";
					when "0010" => out3<= "11011010"; 
					when "0011" => out3<= "11110010"; 
					when "0100" => out3<= "01100110"; 
					when "0101" => out3<= "10110110";
					when "0110" => out3<= "10111110";
					when "0111" => out3<= "11100000"; 
					when "1000" => out3<= "11111110";
					when "1001" => out3<= "11110110";
					when others =>out3<= "01100000";
				end case;
			end if;
		end if;
	end process;
end behavior;